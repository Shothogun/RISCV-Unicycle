package reg_pkg is

type Reg is array (0 to 31)  of bit_vector(31 downto 0);

end reg_pkg;